// injected_biases.vh
localparam logic signed [1*8-1:0] INJECTED_BIASES = 8'sh00;