// injected_weights.vh
localparam logic signed [1*1*2-1:0] INJECTED_WEIGHTS = 2'sh1;